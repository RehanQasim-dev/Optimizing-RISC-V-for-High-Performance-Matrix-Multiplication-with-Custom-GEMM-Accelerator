`timescale 1ns/1ns
module inst_mem_tb;
	logic [31:0] instruction, out;
	
	inst_mem UUT(instruction,out);
		initial begin 
			instruction = 31'h0000_0000;
			#1;
			instruction = 31'h0000_0004;
			#1;
			instruction = 31'h0000_0008;
			#1;
			instruction = 31'h0000_000c;
			#1;
			instruction = 31'h0000_0010;
			#1;
			instruction = 31'h0000_0014;
			#1;
			instruction = 31'h0000_0018;
			#1;
			instruction = 31'h0000_001c;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			instruction = instruction+32'd4;
			#1;
			
			$stop;

		end
endmodule 